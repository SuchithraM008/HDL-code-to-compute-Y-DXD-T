module Test_Bench_DXDT;
parameter N = 8;
reg clk,reset,rst;
reg [7:0]Count;
wire done;
reg [N-1:0]X[63:0];
wire [N+11:0]Y00,Y01,Y02,Y03,Y04,Y05,Y06,Y07,Y10,Y11,Y12,Y13,Y14,Y15,Y16,Y17,Y20,Y21,Y22,Y23,Y24,Y25,Y26,Y27,Y30,Y31,Y32,Y33,Y34,Y35,Y36,Y37,Y40,Y41,Y42,Y43,Y44,Y45,Y46,Y47,Y50,Y51,Y52,Y53,Y54,Y55,Y56,Y57,Y60,Y61,Y62,Y63,Y64,Y65,Y66,Y67,Y70,Y71,Y72,Y73,Y74,Y75,Y76,Y77;

DXDT #(.N(N)) Call_1 (.X00(X[0]),.X01(X[1]),.X02(X[2]),.X03(X[3]),.X04(X[4]),.X05(X[5]),.X06(X[6]),.X07(X[7]),.X10(X[8]),.X11(X[9]),.X12(X[10]),.X13(X[11]),.X14(X[12]),.X15(X[13]),.X16(X[14]),.X17(X[15]),.X20(X[16]),.X21(X[17]),.X22(X[18]),.X23(X[19]),.X24(X[20]),.X25(X[21]),.X26(X[22]),.X27(X[23]),.X30(X[24]),.X31(X[25]),.X32(X[26]),.X33(X[27]),.X34(X[28]),.X35(X[29]),.X36(X[30]),.X37(X[31]),.X40(X[32]),.X41(X[33]),.X42(X[34]),.X43(X[35]),.X44(X[36]),.X45(X[37]),.X46(X[38]),.X47(X[39]),.X50(X[40]),.X51(X[41]),.X52(X[42]),.X53(X[43]),.X54(X[44]),.X55(X[45]),.X56(X[46]),.X57(X[47]),.X60(X[48]),.X61(X[49]),.X62(X[50]),.X63(X[51]),.X64(X[52]),.X65(X[53]),.X66(X[54]),.X67(X[55]),.X70(X[56]),.X71(X[57]),.X72(X[58]),.X73(X[59]),.X74(X[60]),.X75(X[61]),.X76(X[62]),.X77(X[63]),.clk(clk),.reset(reset),.done(done),.Y00(Y00),.Y01(Y01),.Y02(Y02),.Y03(Y03),.Y04(Y04),.Y05(Y05),.Y06(Y06),.Y07(Y07),.Y10(Y10),.Y11(Y11),.Y12(Y12),.Y13(Y13),.Y14(Y14),.Y15(Y15),.Y16(Y16),.Y17(Y17),.Y20(Y20),.Y21(Y21),.Y22(Y22),.Y23(Y23),.Y24(Y24),.Y25(Y25),.Y26(Y26),.Y27(Y27),.Y30(Y30),.Y31(Y31),.Y32(Y32),.Y33(Y33),.Y34(Y34),.Y35(Y35),.Y36(Y36),.Y37(Y37),.Y40(Y40),.Y41(Y41),.Y42(Y42),.Y43(Y43),.Y44(Y44),.Y45(Y45),.Y46(Y46),.Y47(Y47),.Y50(Y50),.Y51(Y51),.Y52(Y52),.Y53(Y53),.Y54(Y54),.Y55(Y55),.Y56(Y56),.Y57(Y57),.Y60(Y60),.Y61(Y61),.Y62(Y62),.Y63(Y63),.Y64(Y64),.Y65(Y65),.Y66(Y66),.Y67(Y67),.Y70(Y70),.Y71(Y71),.Y72(Y72),.Y73(Y73),.Y74(Y74),.Y75(Y75),.Y76(Y76),.Y77(Y77));

initial
begin
clk=1'b1;
repeat(4)
begin
rst=1'b1;
#2700;
end
$stop;
end
always @(posedge clk)
begin
if(rst==1'b1)
begin
Count=8'd0;
reset=1'b1;
rst=1'b0;
end
else if(Count<64)
begin
X[Count]=$random%8;
Count=Count+1'b1;
end
else if(Count==64)
reset=1'b0;
end
always
#5 clk=~clk;

endmodule





           
   
                        